module dc7 (q, d);
output [6:0] q;
input [3:0] d;
assign q[0] = (~d[3] & ~d[2] & ~d[1] & d[0])|(~d[3] & d[2] & ~d[1] &~d[0]); // сегмент а
assign q[1] = (~d[3] & d[2] & ~d[1] & d[0])|(~d[3] & d[2] & d[1] & ~d[0]); // сегмент b
assign q[2] = (~d[3] & ~d[2] & d[1] & ~d[0]); // сегмент c
assign q[3] = (~d[3] & ~d[2] & ~d[1] & d[0])|(~d[3] & d[2] & ~d[1] & ~d[0])|(~d[3] &d[2] & d[1] & d[0]); // сегмент d
assign q[4] = (~d[3] & d[0])|(~d[3] & d[2] & ~d[1])|(~d[2] & ~d[1] & d[0]); // сегмент e
assign q[5] = (~d[3] & ~d[2] & d[0])|(~d[3] & ~d[2] & d[1])|(~d[3] & d[1] & d[0]); //сегмент f
assign q[6] = (~d[3] & ~d[2] & ~d[1])|(~d[3] & d[2] & d[1] & d[0]); // сегмент g
endmodule