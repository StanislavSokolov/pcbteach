-- simple_struct.vhd

-- Generated using ACDS version 22.1 915

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity simple_struct is
	port (
		buzz_buzz             : out std_logic;                                       --       buzz.buzz
		clk_clk               : in  std_logic                    := '0';             --        clk.clk
		enable_enable         : in  std_logic_vector(3 downto 0) := (others => '0'); --     enable.enable
		indicator_indicator   : out std_logic_vector(3 downto 0);                    --  indicator.indicator
		indicator3_indicator3 : in  std_logic_vector(7 downto 0) := (others => '0'); -- indicator3.indicator3
		input0_input0         : in  std_logic                    := '0';             --     input0.input0
		input0_1_input0       : in  std_logic                    := '0';             --   input0_1.input0
		leds_leds             : out std_logic_vector(3 downto 0);                    --       leds.leds
		reset_reset_n         : in  std_logic                    := '0';             --      reset.reset_n
		scl_in                : in  std_logic                    := '0';             --        scl.in
		scl_oe                : out std_logic;                                       --           .oe
		sda_in                : in  std_logic                    := '0';             --        sda.in
		sda_oe                : out std_logic;                                       --           .oe
		segment_segment       : out std_logic_vector(7 downto 0);                    --    segment.segment
		usart_rxd             : in  std_logic                    := '0';             --      usart.rxd
		usart_txd             : out std_logic                                        --           .txd
	);
end entity simple_struct;

architecture rtl of simple_struct is
	component Count250000 is
		port (
			clkIn  : in  std_logic := 'X'; -- clk
			clkOut : out std_logic         -- clk
		);
	end component Count250000;

	component DataConversionUnit is
		port (
			clk        : in  std_logic                    := 'X';             -- clk
			data       : in  std_logic_vector(7 downto 0) := (others => 'X'); -- data
			indicator0 : out std_logic_vector(7 downto 0);                    -- indic0
			indicator1 : out std_logic_vector(7 downto 0);                    -- indic1
			update     : in  std_logic                    := 'X';             -- clk
			indicator2 : out std_logic_vector(7 downto 0)                     -- indic2
		);
	end component DataConversionUnit;

	component DigitalFilter is
		generic (
			PHASE_SHIFT : integer := 2000
		);
		port (
			clk     : in  std_logic := 'X'; -- clk
			output0 : out std_logic;        -- key
			input0  : in  std_logic := 'X'  -- input0
		);
	end component DigitalFilter;

	component DynamicIllumination4Indicators is
		port (
			indicator  : out std_logic_vector(3 downto 0);                    -- indicator
			enable     : in  std_logic_vector(3 downto 0) := (others => 'X'); -- enable
			indicator0 : in  std_logic_vector(7 downto 0) := (others => 'X'); -- indic0
			indicator1 : in  std_logic_vector(7 downto 0) := (others => 'X'); -- indic1
			indicator2 : in  std_logic_vector(7 downto 0) := (others => 'X'); -- indic2
			indicator3 : in  std_logic_vector(7 downto 0) := (others => 'X'); -- indicator3
			segment    : out std_logic_vector(7 downto 0);                    -- segment
			clk        : in  std_logic                    := 'X'              -- clk
		);
	end component DynamicIllumination4Indicators;

	component controller is
		port (
			clk           : in    std_logic                     := 'X';             -- clk
			en            : in    std_logic                     := 'X';             -- reset_n
			uart_rx_busy  : in    std_logic                     := 'X';             -- rx_busy
			uart_rx_data  : in    std_logic_vector(15 downto 0) := (others => 'X'); -- rx_data
			uart_rx_ready : in    std_logic                     := 'X';             -- rx_ready
			uart_tx_data  : out   std_logic_vector(15 downto 0);                    -- tx_data
			uart_tx_dv    : out   std_logic;                                        -- tx_dv
			uart_tx_ready : in    std_logic                     := 'X';             -- tx_ready
			i2c_ack_error : inout std_logic                     := 'X';             -- ack_error
			i2c_addr      : out   std_logic_vector(6 downto 0);                     -- addr
			i2c_busy      : in    std_logic                     := 'X';             -- busy
			i2c_data_rd   : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- data_rd
			i2c_data_wr   : out   std_logic_vector(7 downto 0);                     -- data_wr
			i2c_ena       : out   std_logic;                                        -- ena
			i2c_rw        : out   std_logic;                                        -- rw
			leds          : out   std_logic_vector(3 downto 0);                     -- leds
			dataToUpdate  : out   std_logic_vector(7 downto 0);                     -- data
			key1          : in    std_logic                     := 'X';             -- key
			key2          : in    std_logic                     := 'X';             -- key
			buzz          : out   std_logic                                         -- buzz
		);
	end component controller;

	component i2c_master is
		generic (
			input_clk : integer := 50000000;
			bus_clk   : integer := 100000
		);
		port (
			clk       : in    std_logic                    := 'X';             -- clk
			reset_n   : in    std_logic                    := 'X';             -- reset_n
			ena       : in    std_logic                    := 'X';             -- ena
			addr      : in    std_logic_vector(6 downto 0) := (others => 'X'); -- addr
			rw        : in    std_logic                    := 'X';             -- rw
			data_wr   : in    std_logic_vector(7 downto 0) := (others => 'X'); -- data_wr
			busy      : out   std_logic;                                       -- busy
			data_rd   : out   std_logic_vector(7 downto 0);                    -- data_rd
			ack_error : inout std_logic                    := 'X';             -- ack_error
			scl_in    : in    std_logic                    := 'X';             -- in
			scl_oe    : out   std_logic;                                       -- oe
			sda_in    : in    std_logic                    := 'X';             -- in
			sda_oe    : out   std_logic                                        -- oe
		);
	end component i2c_master;

	component usart is
		generic (
			CLK_FREQ_HZ : integer := 50000000;
			BAUD_RATE   : integer := 9600;
			DATA_BITS   : integer := 8;
			PARITY      : integer := 0;
			STOP_BITS   : integer := 1
		);
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			rx       : in  std_logic                     := 'X';             -- rxd
			tx       : out std_logic;                                        -- txd
			tx_data  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- tx_data
			rx_data  : out std_logic_vector(15 downto 0);                    -- rx_data
			tx_dv    : in  std_logic                     := 'X';             -- tx_dv
			rx_dv    : out std_logic;                                        -- rx_ready
			rx_busy  : out std_logic;                                        -- rx_busy
			tx_ready : out std_logic;                                        -- tx_ready
			en       : in  std_logic                     := 'X'              -- reset_n
		);
	end component usart;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal count250000_0_clkout_clk                 : std_logic;                     -- Count250000_0:clkOut -> DataConversionUnit_0:update
	signal controller_0_datatoupdate_data           : std_logic_vector(7 downto 0);  -- controller_0:dataToUpdate -> DataConversionUnit_0:data
	signal dataconversionunit_0_indic0_indic0       : std_logic_vector(7 downto 0);  -- DataConversionUnit_0:indicator0 -> DynamicIllumination4Indicators_0:indicator0
	signal dataconversionunit_0_indic1_indic1       : std_logic_vector(7 downto 0);  -- DataConversionUnit_0:indicator1 -> DynamicIllumination4Indicators_0:indicator1
	signal dataconversionunit_0_indic2_indic2       : std_logic_vector(7 downto 0);  -- DataConversionUnit_0:indicator2 -> DynamicIllumination4Indicators_0:indicator2
	signal digitalfilter_0_output0_key              : std_logic;                     -- DigitalFilter_0:output0 -> controller_0:key1
	signal digitalfilter_1_output0_key              : std_logic;                     -- DigitalFilter_1:output0 -> controller_0:key2
	signal i2c_transcever_0_port_data_rd            : std_logic_vector(7 downto 0);  -- i2c_transcever_0:data_rd -> controller_0:i2c_data_rd
	signal controller_0_i2c_port_rw                 : std_logic;                     -- controller_0:i2c_rw -> i2c_transcever_0:rw
	signal controller_0_i2c_port_data_wr            : std_logic_vector(7 downto 0);  -- controller_0:i2c_data_wr -> i2c_transcever_0:data_wr
	signal i2c_transcever_0_port_busy               : std_logic;                     -- i2c_transcever_0:busy -> controller_0:i2c_busy
	signal controller_0_i2c_port_ena                : std_logic;                     -- controller_0:i2c_ena -> i2c_transcever_0:ena
	signal controller_0_i2c_port_addr               : std_logic_vector(6 downto 0);  -- controller_0:i2c_addr -> i2c_transcever_0:addr
	signal controller_0_i2c_port_ack_error          : std_logic;                     -- [] -> [controller_0:i2c_ack_error, i2c_transcever_0:ack_error]
	signal usart_0_usart_port_rx_data               : std_logic_vector(15 downto 0); -- usart_0:rx_data -> controller_0:uart_rx_data
	signal usart_0_usart_port_rx_busy               : std_logic;                     -- usart_0:rx_busy -> controller_0:uart_rx_busy
	signal controller_0_uart_port_tx_data           : std_logic_vector(15 downto 0); -- controller_0:uart_tx_data -> usart_0:tx_data
	signal controller_0_uart_port_tx_dv             : std_logic;                     -- controller_0:uart_tx_dv -> usart_0:tx_dv
	signal usart_0_usart_port_rx_ready              : std_logic;                     -- usart_0:rx_dv -> controller_0:uart_rx_ready
	signal usart_0_usart_port_tx_ready              : std_logic;                     -- usart_0:tx_ready -> controller_0:uart_tx_ready
	signal rst_controller_reset_out_reset           : std_logic;                     -- rst_controller:reset_out -> rst_controller_reset_out_reset:in
	signal reset_reset_n_ports_inv                  : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal rst_controller_reset_out_reset_ports_inv : std_logic;                     -- rst_controller_reset_out_reset:inv -> [controller_0:en, i2c_transcever_0:reset_n, usart_0:en]

begin

	count250000_0 : component Count250000
		port map (
			clkIn  => clk_clk,                  --  clkIn.clk
			clkOut => count250000_0_clkout_clk  -- clkOut.clk
		);

	dataconversionunit_0 : component DataConversionUnit
		port map (
			clk        => clk_clk,                            --  clock.clk
			data       => controller_0_datatoupdate_data,     --   data.data
			indicator0 => dataconversionunit_0_indic0_indic0, -- indic0.indic0
			indicator1 => dataconversionunit_0_indic1_indic1, -- indic1.indic1
			update     => count250000_0_clkout_clk,           -- update.clk
			indicator2 => dataconversionunit_0_indic2_indic2  -- indic2.indic2
		);

	digitalfilter_0 : component DigitalFilter
		generic map (
			PHASE_SHIFT => 200
		)
		port map (
			clk     => clk_clk,                     --   clock.clk
			output0 => digitalfilter_0_output0_key, -- output0.key
			input0  => input0_input0                --  input0.input0
		);

	digitalfilter_1 : component DigitalFilter
		generic map (
			PHASE_SHIFT => 2000
		)
		port map (
			clk     => clk_clk,                     --   clock.clk
			output0 => digitalfilter_1_output0_key, -- output0.key
			input0  => input0_1_input0              --  input0.input0
		);

	dynamicillumination4indicators_0 : component DynamicIllumination4Indicators
		port map (
			indicator  => indicator_indicator,                --  indicator.indicator
			enable     => enable_enable,                      --     enable.enable
			indicator0 => dataconversionunit_0_indic0_indic0, -- indicator0.indic0
			indicator1 => dataconversionunit_0_indic1_indic1, -- indicator1.indic1
			indicator2 => dataconversionunit_0_indic2_indic2, -- indicator2.indic2
			indicator3 => indicator3_indicator3,              -- indicator3.indicator3
			segment    => segment_segment,                    --    segment.segment
			clk        => clk_clk                             --        clk.clk
		);

	controller_0 : component controller
		port map (
			clk           => clk_clk,                                  --        clock.clk
			en            => rst_controller_reset_out_reset_ports_inv, --      reset_n.reset_n
			uart_rx_busy  => usart_0_usart_port_rx_busy,               --    uart_port.rx_busy
			uart_rx_data  => usart_0_usart_port_rx_data,               --             .rx_data
			uart_rx_ready => usart_0_usart_port_rx_ready,              --             .rx_ready
			uart_tx_data  => controller_0_uart_port_tx_data,           --             .tx_data
			uart_tx_dv    => controller_0_uart_port_tx_dv,             --             .tx_dv
			uart_tx_ready => usart_0_usart_port_tx_ready,              --             .tx_ready
			i2c_ack_error => controller_0_i2c_port_ack_error,          --     i2c_port.ack_error
			i2c_addr      => controller_0_i2c_port_addr,               --             .addr
			i2c_busy      => i2c_transcever_0_port_busy,               --             .busy
			i2c_data_rd   => i2c_transcever_0_port_data_rd,            --             .data_rd
			i2c_data_wr   => controller_0_i2c_port_data_wr,            --             .data_wr
			i2c_ena       => controller_0_i2c_port_ena,                --             .ena
			i2c_rw        => controller_0_i2c_port_rw,                 --             .rw
			leds          => leds_leds,                                --         leds.leds
			dataToUpdate  => controller_0_datatoupdate_data,           -- dataToUpdate.data
			key1          => digitalfilter_0_output0_key,              --         key1.key
			key2          => digitalfilter_1_output0_key,              --         key2.key
			buzz          => buzz_buzz                                 --         buzz.buzz
		);

	i2c_transcever_0 : component i2c_master
		generic map (
			input_clk => 50000000,
			bus_clk   => 100000
		)
		port map (
			clk       => clk_clk,                                  -- clock.clk
			reset_n   => rst_controller_reset_out_reset_ports_inv, -- reset.reset_n
			ena       => controller_0_i2c_port_ena,                --  port.ena
			addr      => controller_0_i2c_port_addr,               --      .addr
			rw        => controller_0_i2c_port_rw,                 --      .rw
			data_wr   => controller_0_i2c_port_data_wr,            --      .data_wr
			busy      => i2c_transcever_0_port_busy,               --      .busy
			data_rd   => i2c_transcever_0_port_data_rd,            --      .data_rd
			ack_error => controller_0_i2c_port_ack_error,          --      .ack_error
			scl_in    => scl_in,                                   --   SCL.in
			scl_oe    => scl_oe,                                   --      .oe
			sda_in    => sda_in,                                   --   SDA.in
			sda_oe    => sda_oe                                    --      .oe
		);

	usart_0 : component usart
		generic map (
			CLK_FREQ_HZ => 50000000,
			BAUD_RATE   => 9600,
			DATA_BITS   => 8,
			PARITY      => 0,
			STOP_BITS   => 1
		)
		port map (
			clk      => clk_clk,                                  --      clock.clk
			rx       => usart_rxd,                                --        ser.rxd
			tx       => usart_txd,                                --           .txd
			tx_data  => controller_0_uart_port_tx_data,           -- usart_port.tx_data
			rx_data  => usart_0_usart_port_rx_data,               --           .rx_data
			tx_dv    => controller_0_uart_port_tx_dv,             --           .tx_dv
			rx_dv    => usart_0_usart_port_rx_ready,              --           .rx_ready
			rx_busy  => usart_0_usart_port_rx_busy,               --           .rx_busy
			tx_ready => usart_0_usart_port_tx_ready,              --           .tx_ready
			en       => rst_controller_reset_out_reset_ports_inv  --      reset.reset_n
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of simple_struct
