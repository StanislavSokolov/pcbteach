library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;

USE work.i2c_pkg.ALL;

entity controller is
	port(
		en			: in  std_logic;
		clk			: in  std_logic;
		leds	 	: out std_logic_vector( 3 downto 0 );
		
		---------- UART signals ----------------
		uart_tx_data 	: out std_logic_vector(15 downto 0); 	-- data for transmittion
		uart_rx_data 	: in  std_logic_vector(15 downto 0); 	-- external data received
		uart_tx_dv		: out std_logic;						-- tx data valid data latched by rising edge
		uart_rx_ready	: in  std_logic;						-- rx data ready, data set by rising edge
		uart_rx_busy	: in  std_logic;						-- rx busy = 1 while reception in progress
		uart_tx_ready 	: in  std_logic;						-- ready for new operation;	
		
		--------- I2C signals ------------------
		i2c_ena       : out     STD_LOGIC;                    --latch in command
		i2c_addr      : out     STD_LOGIC_VECTOR(6 DOWNTO 0); --address of target slave
		i2c_rw        : out     STD_LOGIC;                    --'0' is write, '1' is read
		i2c_data_wr   : out     STD_LOGIC_VECTOR(7 DOWNTO 0); --data to write to slave
		i2c_busy      : in    	STD_LOGIC;                    --indicates transaction in progress
		i2c_data_rd   : in    	STD_LOGIC_VECTOR(7 DOWNTO 0); --data read from slave
		i2c_ack_error : inout	STD_LOGIC;                    --flag if improper acknowledge from slave
		
		key1 : in STD_LOGIC;									--start
		key2 : in STD_LOGIC;									--stop
		
		dataToUpdate : out STD_LOGIC_VECTOR(7 DOWNTO 0);
		
		buzz : out std_logic
		
	);
end controller;

	
architecture behave of controller is

	CONSTANT CLK_FREQ_HZ 		: INTEGER := 50_000_000;
	CONSTANT UART_BAUDRATE		: INTEGER := 9600;
	constant CLK_I2C_HZ			: INTEGER := 100_000;
	
	CONSTANT wait_500ms  		: INTEGER := CLK_FREQ_HZ / 2;  
	--CONSTANT wait_5ms			: INTEGER := CLK_FREQ_HZ / 200;
	
	CONSTANT wait_05ms  		: INTEGER := CLK_FREQ_HZ / 25000; -- 1000 Hz
	CONSTANT wait_1ms  		: INTEGER := CLK_FREQ_HZ / 50000; -- 500 Hz
	
	constant I2C_SLAVE_ADDR 	: STD_LOGIC_VECTOR( 6 DOWNTO 0 ) := "1001000";
	constant TEMPER_REG_ADDR	: STD_LOGIC_VECTOR( 7 DOWNTO 0 ) := x"00";
	
	
	
	component pgen IS		-- 1 cicle pulse generator
	GENERIC(
		Edge : STD_LOGIC	-- 0 = falling edge, 1 = rising edge pulse gen
	);
	PORT(
		Enable : IN  STD_LOGIC;
		Clk    : IN  STD_LOGIC;
		Input  : IN  STD_LOGIC;
		Output : OUT STD_LOGIC
	);
	END component pgen;
	
	
	
	

		
		
	SIGNAL wait_cnt				: integer range 0 to wait_500ms;
	SIGNAL tx_start				: std_logic;
	SIGNAL dv_cnt 				: integer range 0 to 2;
	SIGNAL symbol_counter  		: integer range 0 to 3;
	
--	signal cnt_100Hz   			: integer range 0 to wait_5ms;
--	signal clk_100Hz			: std_logic;
--	signal btn_cnt              : integer range 0 to 4;

	signal cnt_500Hz   			: integer range 0 to wait_1ms;
	signal clk_500Hz			: std_logic;
	
	signal cnt_1000Hz   			: integer range 0 to wait_05ms;
	signal clk_1000Hz			: std_logic;

	signal cnt_05Hz   			: integer range 0 to CLK_FREQ_HZ;
	signal clk_05Hz			: std_logic;	
	
	type FSM_State	is 	( IDLE, READ_TEMPER, UPDATE_IND, SEND_TEMPER, SEND_LIMIT );
	signal PresState : FSM_State;
	
	signal reset_n   :   STD_LOGIC;                    --active low reset

	signal count_1Hz 	: integer range 0 to wait_500ms;
	signal clk_1Hz		: STD_LOGIC;
	signal StartPulse	: STD_LOGIC;
	
	
	signal sda_line		: STD_LOGIC;
	signal scl_line		: STD_LOGIC;
	
	SIGNAL I2C_RxDataLen : INTEGER RANGE 0 TO I2C_DATA_LEN_MAX;
	SIGNAL I2C_RxArray   : I2C_Rd_Array;
	SIGNAL RxByteCnt     : INTEGER RANGE 0 TO 15;
	
	SIGNAL I2C_ByteCnt : INTEGER RANGE 0 TO I2C_DATA_LEN_MAX;
	SIGNAL I2C_PackLen : INTEGER RANGE 0 TO 63;
	
	SIGNAL RegWrDone 	: STD_LOGIC;
	SIGNAL RegRdDone 	: STD_LOGIC;
	SIGNAL I2C_BusyPrev : STD_LOGIC;
	
	
	SIGNAL I2C_Load      : STD_LOGIC;
	signal I2C_DevAddr  : STD_LOGIC_VECTOR( I2C_ADDR_WIDTH-1 DOWNTO 0 );	
	signal I2C_WrData   : STD_LOGIC_VECTOR( I2C_DATA_WIDTH-1 DOWNTO 0 );	
	signal I2C_RdData   : STD_LOGIC_VECTOR( I2C_DATA_WIDTH-1 DOWNTO 0 );	
	signal I2C_Err      : STD_LOGIC;	
	
	SIGNAL Temper  		: STD_LOGIC_VECTOR( 7 DOWNTO 0 );
	SIGNAL Temper_Limit_Low  		: STD_LOGIC_VECTOR( 7 DOWNTO 0 ) := x"14"; -- 20 градусов
	SIGNAL Temper_Limit_High  		: STD_LOGIC_VECTOR( 7 DOWNTO 0 ) := x"1E"; -- 30 градусов
	SIGNAL CMD : STD_LOGIC_VECTOR( 7 DOWNTO 0 ) := x"F0";
	SIGNAL send_limit_en : STD_LOGIC := '0';
	
	SIGNAL key1Prev : STD_LOGIC := '0';
	SIGNAL key2Prev : STD_LOGIC := '0';
	SIGNAL start_stop : STD_LOGIC := '1';
	
	SIGNAL buzz_mode : STD_LOGIC_VECTOR(1 DOWNTO 0) := b"00";
	
	
	SIGNAL cmdLimit : STD_LOGIC := '0';
	SIGNAL uart_rx_ready_prev : STD_LOGIC := '0';

begin

	 
	
	start_gen: pgen 		-- 1 cicle pulse generator
	GENERIC MAP(
		Edge => '1' 	--  1 = rising edge pulse gen
	)
	PORT MAP(
		Enable 	=>	reset_n	,
		Clk    	=>	clk		,
		Input  	=>	clk_1Hz		,
		Output 	=>	StartPulse		-- generate start pulse 1 cicle clk width every second 
	);
	
		
	reset_n	<= en;
	
	
	i2c_ena     	<=	 I2C_Load    ;
	i2c_addr    	<=	 I2C_DevAddr ;
--	i2c_rw_int      <=	 I2C_RW      ;
	i2c_data_wr 	<=	 I2C_WrData  ;
--	I2C_Busy_int   	<=	i2c_busy      ;
	I2C_RdData 		<=	i2c_data_rd   ;
	I2C_Err    		<=	i2c_ack_error ;
	
	gen_start_stop: process( reset_n, clk )
	begin
		if reset_n = '0' then
			start_stop <= '0';
		elsif rising_edge( clk ) then
			if key1 = '0' and key1Prev = '1' then
				start_stop <= '1';
			elsif key2 = '0' and key2Prev = '1' then
				start_stop <= '0';
			end if;
			key1Prev <= key1;
			key2Prev <= key2;				
		end if;
	end process;	
	
	gen_05Hz: process( reset_n, clk )
	begin
		if reset_n = '0' then
			cnt_05Hz 	<= 0;
			clk_05Hz		<= '0';
		elsif rising_edge( clk ) then
			if cnt_05Hz < CLK_FREQ_HZ then
				cnt_05Hz <= cnt_05Hz + 1;
			else	
				cnt_05Hz <= 0;
				clk_05Hz <= NOT clk_05Hz;
			end if;
		end if;
	end process;

	gen_500Hz: process( reset_n, clk )
	begin
		if reset_n = '0' then
			cnt_500Hz 	<= 0;
			clk_500Hz		<= '0';
		elsif rising_edge( clk ) then
			if cnt_500Hz < wait_1ms then
				cnt_500Hz <= cnt_500Hz + 1;
			else	
				cnt_500Hz <= 0;
				clk_500Hz <= NOT clk_500Hz;
			end if;
		end if;
	end process;

	gen_1000Hz: process( reset_n, clk )
	begin
		if reset_n = '0' then
			cnt_1000Hz 	<= 0;
			clk_1000Hz		<= '0';
		elsif rising_edge( clk ) then
			if cnt_1000Hz < wait_05ms then
				cnt_1000Hz <= cnt_1000Hz + 1;
			else	
				cnt_1000Hz <= 0;
				clk_1000Hz <= NOT clk_1000Hz;
			end if;
		end if;
	end process;	
	
	gen_1Hz: process( reset_n, clk )
	begin
		if reset_n = '0' then
			count_1Hz 	<= 0;
			clk_1Hz		<= '0';
		elsif rising_edge( clk ) then
			if count_1Hz < wait_500ms then
				count_1Hz <= count_1Hz + 1;
			else	
				count_1Hz <= 0;
				clk_1Hz <= NOT clk_1Hz;
			end if;
		end if;
	end process;
	
	work_buzz: process( reset_n, clk )
	begin
		if reset_n = '0' then
			buzz <= '0';
		elsif rising_edge( clk ) then
			case buzz_mode is
				when b"01" =>
					buzz <= clk_05Hz and clk_500Hz;
				when b"10" => 
					buzz <= clk_05Hz and clk_1000Hz; 	
				when others =>
					buzz <= '0';
			end case;				
		end if;
	end process;
	
	ReceiveCMD: process( reset_n, clk )
		variable byteCount : integer range 0 to 1 := 0;
	begin
		if reset_n = '0' then
			byteCount := 0;
		elsif rising_edge( clk ) then
			IF uart_rx_busy = '0' and uart_rx_ready = '1' and uart_rx_ready_prev = '0' THEN 
				if byteCount = 0 then
					cmdLimit <= uart_rx_data(0);
					byteCount := 1;
				else
					if cmdLimit = '0' then
						Temper_Limit_Low <= uart_rx_data(7 downto 0);
					else 
						Temper_Limit_High <= uart_rx_data(7 downto 0);
					end if;
					byteCount := 0;
				end if;		
			end if;
			uart_rx_ready_prev <= uart_rx_ready;
		end if;
	end process;
	

	FSM: process( reset_n, clk )
		variable show_cnt : integer range 0 to 25;
		
	begin
		if reset_n = '0' or start_stop = '0' then
			PresState <= IDLE;
			show_cnt 	:= 0;
			Temper		 <= ( others => '0' );
			buzz_mode <= b"11";
			uart_tx_dv 		<= '0';
		elsif rising_edge( clk ) then
		
			I2C_BusyPrev <= I2C_Busy;
			
			case ( PresState ) is
			
			when IDLE =>
				I2C_Load 	<= '0';
				I2C_ByteCnt <= 0;
				RegWrDone  	<= '0';
				RegRdDone  	<= '0';
				I2C_BusyPrev <= '0';
				
				show_cnt 	:= 0;
				
				I2C_RxDataLen <= 2;
				
				uart_tx_dv 		<= '0';	

				
	
				IF uart_tx_ready = '1' THEN
					IF send_limit_en = '1' THEN
						send_limit_en <= '0';
						IF Temper_Limit_Low <= Temper_Limit_High THEN
							IF Temper < Temper_Limit_Low THEN
								CMD <= x"F1";							-- превышен нижний порог
								leds <= b"1110";
								buzz_mode <= b"01";
							ELSE 
								IF Temper >	Temper_Limit_High THEN
									CMD <= x"F2";						-- превышен верхний порог
									leds <= b"0111";
									buzz_mode <= b"10";
								ELSE
									CMD <= x"F0";						-- темпреатура в норме
									leds <= b"1001";
									buzz_mode <= b"00";
								END IF;
							END IF;
						ELSE
							CMD <= x"F3";								-- неверно заданы пределы температуры
						END IF;									
						PresState <= SEND_LIMIT;
					ELSE	
						IF I2C_Busy = '0' THEN
							IF StartPulse = '1' THEN
								PresState <= READ_TEMPER; 
							END IF;
						END IF;
					END IF;		
				END IF;
			
			when READ_TEMPER =>
				if RegRdDone = '0' then    
					i2c_array_rd( 
				          I2C_SLAVE_ADDR,    -- I2C Bus device Address
	                      TEMPER_REG_ADDR, -- I2C device internal register address
	                      I2C_RxArray,		   -- I2C device temper readed 2 bytes
	                      I2C_ByteCnt,          -- Byte Counter
						  I2C_RxDataLen,		-- Rx Array len = 2 bytes
	                      I2C_DevAddr,         
	                      I2C_RW,              
	                      I2C_Load,             
	                      I2C_Busy,            
	                      I2C_BusyPrev,        
	                      RegRdDone,           -- Data Read Ready Flag
	                      I2C_WrData,
	                      I2C_RdData           
	                );
					PresState <= READ_TEMPER;
				
				elsif I2C_Err = '0' then
					Temper 		<= I2C_RxArray(0);	-- use MSB of readed temper value. It's in integer temper value
					RegRdDone 	<= '0';
					PresState 	<= UPDATE_IND;
				else
					PresState <= IDLE;
					
				end if;
				
			when UPDATE_IND =>
				dataToUpdate <= Temper;
				PresState 	<= SEND_TEMPER;
			
			when SEND_TEMPER =>
				if show_cnt < 2 then
					show_cnt := show_cnt + 1;
					
					uart_tx_dv 		<= '1';
					uart_tx_data( 7 downto 0 ) 	<= Temper;
					PresState 		<= SEND_TEMPER;
				else
					uart_tx_dv 		<= '0';
					show_cnt := 0;
					PresState <= IDLE;
					send_limit_en <= '1';
				end if;
				
			when SEND_LIMIT =>
				if show_cnt < 2 then
					show_cnt := show_cnt + 1;
					
					uart_tx_dv 		<= '1';
					uart_tx_data( 7 downto 0 ) 	<= CMD;
					PresState 		<= SEND_LIMIT;
				else
					uart_tx_dv 		<= '0';
					show_cnt := 0;
					PresState <= IDLE;
				end if;	
			
			when OTHERS => 
				PresState <= IDLE;
				
			end case;
			
		
		end if;
	
	
	end process;
	
	
	
	
	
	
end behave;