LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY IPblock IS 
	PORT
	(
		clk :  IN  STD_LOGIC;
		key1 :  IN  STD_LOGIC;
		key2 :  IN  STD_LOGIC;
		led1 :  OUT  STD_LOGIC;
		led2 :  OUT  STD_LOGIC;
		led3 :  OUT  STD_LOGIC;
		buzz :  OUT  STD_LOGIC
	);
END IPblock;

ARCHITECTURE bdf_type OF IPblock IS 

COMPONENT altpll01
	PORT(inclk0 : IN STD_LOGIC;
		 areset : IN STD_LOGIC;
		 c0 : OUT STD_LOGIC;
		 locked : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT dtrigwre
	PORT(D : IN STD_LOGIC;
		 C : IN STD_LOGIC;
		 Q : OUT STD_LOGIC;
		 nQ : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT countm1
	PORT(clock : IN STD_LOGIC;
		 cout : OUT STD_LOGIC;
		 q : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END COMPONENT;

COMPONENT countm9
	PORT(clock : IN STD_LOGIC;
		 cout : OUT STD_LOGIC;
		 q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	);
END COMPONENT;

COMPONENT logblock
	PORT(clk : IN STD_LOGIC;
		 input0 : IN STD_LOGIC;
		 input1 : IN STD_LOGIC;
		 output : OUT STD_LOGIC
	);
END COMPONENT;

COMPONENT countm2
	PORT(clock : IN STD_LOGIC;
		 cout : OUT STD_LOGIC;
		 q : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	SYNTHESIZED_WIRE_0 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;


BEGIN 
SYNTHESIZED_WIRE_0 <= '0';



b2v_inst : altpll01
PORT MAP(inclk0 => clk,
		 areset => SYNTHESIZED_WIRE_0,
		 c0 => SYNTHESIZED_WIRE_10);


b2v_inst1 : dtrigwre
PORT MAP(D => SYNTHESIZED_WIRE_1,
		 C => SYNTHESIZED_WIRE_20,
		 Q => SYNTHESIZED_WIRE_7,
		 nQ => SYNTHESIZED_WIRE_1);


b2v_inst10 : countm1
PORT MAP(clock => SYNTHESIZED_WIRE_21,
		 cout => SYNTHESIZED_WIRE_19);


b2v_inst11 : dtrigwre
PORT MAP(D => SYNTHESIZED_WIRE_4,
		 C => SYNTHESIZED_WIRE_21,
		 Q => led3,
		 nQ => SYNTHESIZED_WIRE_4);


buzz <= SYNTHESIZED_WIRE_6 AND SYNTHESIZED_WIRE_7;


b2v_inst14 : dtrigwre
PORT MAP(D => SYNTHESIZED_WIRE_8,
		 C => key1,
		 Q => SYNTHESIZED_WIRE_13,
		 nQ => SYNTHESIZED_WIRE_8);


b2v_inst15 : dtrigwre
PORT MAP(D => SYNTHESIZED_WIRE_9,
		 C => key2,
		 Q => SYNTHESIZED_WIRE_14,
		 nQ => SYNTHESIZED_WIRE_9);



b2v_inst3 : countm9
PORT MAP(clock => SYNTHESIZED_WIRE_10,
		 cout => SYNTHESIZED_WIRE_20);


b2v_inst4 : countm9
PORT MAP(clock => SYNTHESIZED_WIRE_20,
		 cout => SYNTHESIZED_WIRE_12);


b2v_inst5 : countm9
PORT MAP(clock => SYNTHESIZED_WIRE_12,
		 cout => SYNTHESIZED_WIRE_21);


b2v_inst6 : logblock
PORT MAP(clk => clk,
		 input0 => SYNTHESIZED_WIRE_13,
		 input1 => SYNTHESIZED_WIRE_14,
		 output => SYNTHESIZED_WIRE_6);


b2v_inst7 : dtrigwre
PORT MAP(D => SYNTHESIZED_WIRE_15,
		 C => SYNTHESIZED_WIRE_16,
		 Q => led1,
		 nQ => SYNTHESIZED_WIRE_15);


b2v_inst8 : countm2
PORT MAP(clock => SYNTHESIZED_WIRE_21,
		 cout => SYNTHESIZED_WIRE_16);


b2v_inst9 : dtrigwre
PORT MAP(D => SYNTHESIZED_WIRE_18,
		 C => SYNTHESIZED_WIRE_19,
		 Q => led2,
		 nQ => SYNTHESIZED_WIRE_18);


END bdf_type;